/*
 This file is top level of Gated Recurrent Unit (GRU).
 This is the part of DLPR32 processor 

*/
module gruMain();
 
  
endmodule
