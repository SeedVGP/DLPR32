/* Floating Point Processor of 16 Bits along with 32bit RISC V*/


module riscvfzfh ();
  input
  output
  
  
  
endmodule
