`timescale 1ns/1ps 
module addss(
input clk,cs_add,rst,
  input [15:0]x,y,
output reg [15:0] sum,
output reg rdy_add
);
reg cout;
reg [15:0] op1,op2;
reg [15:0] p,g,c;
reg [1:0] state=0;

always@(posedge clk)
begin
if(rst)
begin
state=0;

end
else
begin
case(state)
0:begin
	if(cs_add)
	state=1;
  	else
	state=0;
  end
1:state=2;
2:state=3;
3:begin
	if(rdy_add)
	state=0;
	else
	state=3;
  end
endcase
end
end
  
always@(state)
begin
case(state)
0:rdy_add=1;
1:rdy_add=0;
2:
  begin
    sum=16'b0;

    op1=x;
    op2=y;
    if(x[15]==1'b1)
      op1={1'b1,~x[14:0]+1'b1};
    else
	op1=op1;
    if(y[15]==1'b1)
      op2={1'b1,~y[14:0]+1'b1};
    else
	op2=op2;
  end
3:begin
 p=op1^op2;
 g=op1&op2;
  c[0]=1'b0;
          
 c[1]=g[0]|(p[0]&c[0]);
          
 c[2]=g[1]|(p[1]&g[0])|(p[1]&p[0]&c[0]);
          
 c[3]=g[2]|(p[2]&g[1])|(p[2]&p[1]&g[0])|(p[2]&p[1]&p[0]&c[0]);
          
 c[4]=g[3]|(p[3]&g[2])|(p[3]&p[2]&g[1])|(p[3]&p[2]&p[1]&g[0])|(p[3]&p[2]&p[1]&p[0]&c[0]);
 
 c[5]=g[4] | (p[4]&g[3]) | (p[4]&p[3]&g[2]) | (p[4]&p[3]&p[2]&g[1]) |(p[4]&p[3]&p[2]&p[1]&g[0]) | (p[4]&p[3]&p[2]&p[1]&p[0]&c[0]); 
          
 c[6]=g[5] | (p[5]&g[4]) | (p[5]&p[4]&g[3]) | (p[5]&p[4]&p[3]&g[2]) | (p[5]&p[4]&p[3]&p[2]&g[1]) | (p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);

 c[7]=g[6] | (p[6]&g[5]) | (p[6]&p[5]&g[4]) | (p[6]&p[5]&p[4]&g[3]) | (p[6]&p[5]&p[4]&p[3]&g[2]) | (p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);

c[8]=g[7] | (p[7]&g[6]) | (p[7]&p[6]&g[5]) | (p[7]&p[6]&p[5]&g[4]) | (p[7]&p[6]&p[5]&p[4]&g[3]) | (p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);

c[9]=g[8] | (p[8]&g[7]) | (p[8]&p[7]&g[6]) | (p[8]&p[7]&p[6]&g[5]) | (p[8]&p[7]&p[6]&p[5]&g[4]) | (p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);

c[10]=g[9] | (p[9]&g[8]) | (p[9]&p[8]&g[7]) | (p[9]&p[8]&p[7]&g[6]) | (p[9]&p[8]&p[7]&p[6]&g[5]) | (p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);

c[11]=g[10] | (p[10]&g[9]) | (p[10]&p[9]&g[8]) | (p[10]&p[9]&p[8]&g[7]) | (p[10]&p[9]&p[8]&p[7]&g[6]) | (p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);
c[12]=g[11] | (p[11]&g[10]) |(p[11]&p[10]&g[9]) | (p[11]&p[10]&p[9]&g[8]) | (p[11]&p[10]&p[9]&p[8]&g[7]) | (p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);
 c[13]=g[12] | (p[12]&g[11]) | (p[12]&p[11]&g[10]) |( p[12]&p[11]&p[10]&g[9]) | (p[12]&p[11]&p[10]&p[9]&g[8]) | (p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);
c[14]=g[13] | (p[13]&g[12]) | (p[13]&p[12]&g[11]) | (p[13]&p[12]&p[11]&g[10]) |( p[13]&p[12]&p[11]&p[10]&g[9]) | (p[13]&p[12]&p[11]&p[10]&p[9]&g[8]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);
c[15]=g[14] | (p[14]&g[13]) |  (p[14]&p[13]&g[12]) | (p[14]&p[13]&p[12]&g[11]) | (p[14]&p[13]&p[12]&p[11]&g[10]) |( p[14]&p[13]&p[12]&p[11]&p[10]&g[9]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);
cout=g[15] | (p[15]&g[14]) | (p[15]&p[14]&g[13]) |  (p[15]&p[14]&p[13]&g[12]) | (p[15]&p[14]&p[13]&p[12]&g[11]) | (p[15]&p[14]&p[13]&p[12]&p[11]&g[10]) |( p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c[0]);
 
 sum=p^c;
  if(sum[15]==1'b1)
    sum={1'b1,~sum[14:0]+1'b1};
  else
	sum=sum;
rdy_add=1;

end
endcase
end
endmodule



//-----------------------------------TEST BENCH----------------------------------------------------------
`timescale 1ns/1ps 
module addss_tb(); 

reg clk,cs_add,rst;
  reg [15:0] x,y;
wire [15:0] sum;
wire rdy_add;
  addss u0(clk,cs_add,rst,x,y,sum,rdy_add);
initial
begin
clk=1'b0;
forever #5 clk=~clk;
end
initial
begin
  //$dumpfile("dump.vcd");
//$dumpvars;
rst=1'b1;
cs_add=0;
#10;
rst=1'b0;
cs_add=1;
x=16'b1011010000000000;
y=16'b1000010000000000;

#100;
$finish;
end
endmodule
