/* Main RISC V Core file */ 


module DRISCV(
  
);
  input clk,Din;
  output Dout;
  // Above is general input and output need to define properly 
  
  // Call for control, Memory and ALU modules from here
  
  
endmodule
